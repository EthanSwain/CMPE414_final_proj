module MADcalc #(parameter scale_factor = 'h017C,)();

endmodule